module mux4to1 (
    input wire a,       
    input wire b,       
    input wire c,        
    input wire d,        
    input wire [1:0] sel,
    output wire y       
);
    assign y = (sel == 2'b00) ? a :
               (sel == 2'b01) ? b :
               (sel == 2'b10) ? c :
                                d;   
endmodule
